library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity B_RAM_0 is
	port (
		clk 		: in std_logic;
		we 			: in std_logic;
		fetch		: in std_logic;
		addr_inst 	: in std_logic_vector (29 downto 0);
		addr_data	: in std_logic_vector (29 downto 0);
		data_in 	: in std_logic_vector (7 downto 0);

		inst_out 	: out std_logic_vector (7 downto 0);
		data_out 	: out std_logic_vector (7 downto 0)
	);
end B_RAM_0;

-- 8 kB BRAM
architecture behavioral of B_RAM_0 is

	type ram_type is array (0 to 8192) of std_logic_vector(7 downto 0);
	signal ram : ram_type := (
		0 => x"97",
		1 => x"93",
		2 => x"73",
		3 => x"17",
		4 => x"13",
		5 => x"ef",
		6 => x"6f",
		7 => x"13",
		8 => x"23",
		9 => x"ef",
		10 => x"ef",
		11 => x"ef",
		12 => x"83",
		13 => x"13",
		14 => x"73",
		15 => x"13",
		16 => x"23",
		17 => x"23",
		18 => x"23",
		19 => x"23",
		20 => x"23",
		21 => x"23",
		22 => x"23",
		23 => x"23",
		24 => x"23",
		25 => x"23",
		26 => x"23",
		27 => x"23",
		28 => x"23",
		29 => x"23",
		30 => x"23",
		31 => x"23",
		32 => x"23",
		33 => x"23",
		34 => x"23",
		35 => x"23",
		36 => x"23",
		37 => x"23",
		38 => x"23",
		39 => x"23",
		40 => x"23",
		41 => x"23",
		42 => x"23",
		43 => x"23",
		44 => x"23",
		45 => x"67",
		46 => x"83",
		47 => x"03",
		48 => x"83",
		49 => x"03",
		50 => x"83",
		51 => x"03",
		52 => x"83",
		53 => x"03",
		54 => x"83",
		55 => x"03",
		56 => x"83",
		57 => x"03",
		58 => x"83",
		59 => x"03",
		60 => x"83",
		61 => x"03",
		62 => x"83",
		63 => x"03",
		64 => x"83",
		65 => x"03",
		66 => x"83",
		67 => x"03",
		68 => x"83",
		69 => x"03",
		70 => x"83",
		71 => x"03",
		72 => x"83",
		73 => x"03",
		74 => x"83",
		75 => x"13",
		76 => x"67",
		77 => x"13",
		78 => x"23",
		79 => x"13",
		80 => x"f3",
		81 => x"23",
		82 => x"83",
		83 => x"13",
		84 => x"03",
		85 => x"13",
		86 => x"67",
		87 => x"13",
		88 => x"23",
		89 => x"13",
		90 => x"23",
		91 => x"83",
		92 => x"73",
		93 => x"13",
		94 => x"03",
		95 => x"13",
		96 => x"67",
		97 => x"13",
		98 => x"23",
		99 => x"13",
		100 => x"23",
		101 => x"83",
		102 => x"73",
		103 => x"13",
		104 => x"03",
		105 => x"13",
		106 => x"67",
		107 => x"13",
		108 => x"23",
		109 => x"13",
		110 => x"23",
		111 => x"83",
		112 => x"73",
		113 => x"13",
		114 => x"03",
		115 => x"13",
		116 => x"67",
		117 => x"13",
		118 => x"23",
		119 => x"13",
		120 => x"23",
		121 => x"83",
		122 => x"73",
		123 => x"13",
		124 => x"03",
		125 => x"13",
		126 => x"67",
		127 => x"13",
		128 => x"23",
		129 => x"13",
		130 => x"f3",
		131 => x"23",
		132 => x"83",
		133 => x"13",
		134 => x"03",
		135 => x"13",
		136 => x"67",
		137 => x"13",
		138 => x"23",
		139 => x"23",
		140 => x"13",
		141 => x"13",
		142 => x"ef",
		143 => x"13",
		144 => x"93",
		145 => x"ef",
		146 => x"ef",
		147 => x"13",
		148 => x"6f",
		149 => x"13",
		150 => x"23",
		151 => x"23",
		152 => x"13",
		153 => x"b7",
		154 => x"03",
		155 => x"83",
		156 => x"03",
		157 => x"83",
		158 => x"b7",
		159 => x"13",
		160 => x"33",
		161 => x"93",
		162 => x"b3",
		163 => x"b3",
		164 => x"b3",
		165 => x"93",
		166 => x"13",
		167 => x"93",
		168 => x"23",
		169 => x"23",
		170 => x"13",
		171 => x"ef",
		172 => x"13",
		173 => x"83",
		174 => x"03",
		175 => x"13",
		176 => x"67",
		177 => x"13",
		178 => x"23",
		179 => x"13",
		180 => x"23",
		181 => x"23",
		182 => x"03",
		183 => x"83",
		184 => x"23",
		185 => x"23",
		186 => x"b7",
		187 => x"03",
		188 => x"83",
		189 => x"03",
		190 => x"83",
		191 => x"b7",
		192 => x"13",
		193 => x"33",
		194 => x"93",
		195 => x"b3",
		196 => x"b3",
		197 => x"b3",
		198 => x"93",
		199 => x"13",
		200 => x"93",
		201 => x"23",
		202 => x"23",
		203 => x"13",
		204 => x"03",
		205 => x"13",
		206 => x"67",
		207 => x"13",
		208 => x"23",
		209 => x"23",
		210 => x"13",
		211 => x"13",
		212 => x"ef",
		213 => x"13",
		214 => x"ef",
		215 => x"13",
		216 => x"83",
		217 => x"03",
		218 => x"13",
		219 => x"67",
		220 => x"13",
		221 => x"23",
		222 => x"13",
		223 => x"23",
		224 => x"23",
		225 => x"6f",
		226 => x"83",
		227 => x"03",
		228 => x"b3",
		229 => x"03",
		230 => x"b7",
		231 => x"23",
		232 => x"83",
		233 => x"93",
		234 => x"23",
		235 => x"83",
		236 => x"03",
		237 => x"b3",
		238 => x"83",
		239 => x"e3",
		240 => x"13",
		241 => x"13",
		242 => x"03",
		243 => x"13",
		244 => x"67",
		245 => x"13",
		246 => x"23",
		247 => x"13",
		248 => x"23",
		249 => x"23",
		250 => x"83",
		251 => x"23",
		252 => x"23",
		253 => x"6f",
		254 => x"03",
		255 => x"83",
		256 => x"b3",
		257 => x"a3",
		258 => x"03",
		259 => x"83",
		260 => x"b3",
		261 => x"23",
		262 => x"83",
		263 => x"93",
		264 => x"13",
		265 => x"83",
		266 => x"93",
		267 => x"b3",
		268 => x"23",
		269 => x"83",
		270 => x"93",
		271 => x"23",
		272 => x"83",
		273 => x"e3",
		274 => x"83",
		275 => x"93",
		276 => x"23",
		277 => x"6f",
		278 => x"83",
		279 => x"93",
		280 => x"b3",
		281 => x"03",
		282 => x"b7",
		283 => x"23",
		284 => x"83",
		285 => x"93",
		286 => x"23",
		287 => x"83",
		288 => x"e3",
		289 => x"13",
		290 => x"13",
		291 => x"03",
		292 => x"13",
		293 => x"67",
		294 => x"13",
		295 => x"23",
		296 => x"23",
		297 => x"13",
		298 => x"ef",
		299 => x"23",
		300 => x"03",
		301 => x"b7",
		302 => x"93",
		303 => x"63",
		304 => x"ef",
		305 => x"6f",
		306 => x"13",
		307 => x"ef",
		308 => x"93",
		309 => x"03",
		310 => x"ef",
		311 => x"13",
		312 => x"ef",
		313 => x"13",
		314 => x"6f",
		315 => x"13",
		316 => x"83",
		317 => x"03",
		318 => x"13",
		319 => x"67",
		320 => x"48",
		321 => x"6f",
		322 => x"72",
		323 => x"0a",
		324 => x"54",
		325 => x"21",
		326 => x"55",
		327 => x"70",
		328 => x"65",
		329 => x"63",
		330 => x"65",
		331 => x"75",
		332 => x"20",
		333 => x"0a",
		others => (others => '0')
	);

begin

	process(clk)
	begin
		if (rising_edge(clk)) then
			if (fetch = '1') then
				inst_out <= ram(to_integer(unsigned(addr_inst(12 downto 0))));
			end if;

			if (we = '1') then
				ram(to_integer(unsigned(addr_data(12 downto 0)))) <= data_in;
			end if;
			
			data_out <= ram(to_integer(unsigned(addr_data(12 downto 0))));
		end if;
	end process;

end behavioral ; -- arch

