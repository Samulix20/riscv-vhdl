library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity B_RAM_2 is
	port (
		clk 		: in std_logic;
		we 			: in std_logic;
		fetch		: in std_logic;
		addr_inst 	: in std_logic_vector (29 downto 0);
		addr_data	: in std_logic_vector (29 downto 0);
		data_in 	: in std_logic_vector (7 downto 0);

		inst_out 	: out std_logic_vector (7 downto 0);
		data_out 	: out std_logic_vector (7 downto 0)
	);
end B_RAM_2;

-- 8 kB BRAM
architecture behavioral of B_RAM_2 is

	type ram_type is array (0 to 8192) of std_logic_vector(7 downto 0);
	signal ram : ram_type := (
		0 => x"00",
		1 => x"c0",
		2 => x"50",
		3 => x"00",
		4 => x"41",
		5 => x"00",
		6 => x"00",
		7 => x"c1",
		8 => x"11",
		9 => x"80",
		10 => x"00",
		11 => x"c0",
		12 => x"01",
		13 => x"41",
		14 => x"20",
		15 => x"c1",
		16 => x"31",
		17 => x"41",
		18 => x"51",
		19 => x"61",
		20 => x"71",
		21 => x"81",
		22 => x"91",
		23 => x"a1",
		24 => x"b1",
		25 => x"c1",
		26 => x"d1",
		27 => x"e1",
		28 => x"f1",
		29 => x"01",
		30 => x"11",
		31 => x"21",
		32 => x"31",
		33 => x"41",
		34 => x"51",
		35 => x"61",
		36 => x"71",
		37 => x"81",
		38 => x"91",
		39 => x"a1",
		40 => x"b1",
		41 => x"c1",
		42 => x"d1",
		43 => x"e1",
		44 => x"f1",
		45 => x"00",
		46 => x"01",
		47 => x"41",
		48 => x"81",
		49 => x"c1",
		50 => x"01",
		51 => x"41",
		52 => x"81",
		53 => x"c1",
		54 => x"01",
		55 => x"41",
		56 => x"81",
		57 => x"c1",
		58 => x"01",
		59 => x"41",
		60 => x"81",
		61 => x"c1",
		62 => x"01",
		63 => x"41",
		64 => x"81",
		65 => x"c1",
		66 => x"01",
		67 => x"41",
		68 => x"81",
		69 => x"c1",
		70 => x"01",
		71 => x"41",
		72 => x"81",
		73 => x"c1",
		74 => x"01",
		75 => x"41",
		76 => x"00",
		77 => x"01",
		78 => x"81",
		79 => x"01",
		80 => x"20",
		81 => x"f4",
		82 => x"c4",
		83 => x"07",
		84 => x"c1",
		85 => x"01",
		86 => x"00",
		87 => x"01",
		88 => x"81",
		89 => x"01",
		90 => x"a4",
		91 => x"c4",
		92 => x"47",
		93 => x"00",
		94 => x"c1",
		95 => x"01",
		96 => x"00",
		97 => x"01",
		98 => x"81",
		99 => x"01",
		100 => x"a4",
		101 => x"c4",
		102 => x"47",
		103 => x"00",
		104 => x"c1",
		105 => x"01",
		106 => x"00",
		107 => x"01",
		108 => x"81",
		109 => x"01",
		110 => x"a4",
		111 => x"c4",
		112 => x"07",
		113 => x"00",
		114 => x"c1",
		115 => x"01",
		116 => x"00",
		117 => x"01",
		118 => x"81",
		119 => x"01",
		120 => x"a4",
		121 => x"c4",
		122 => x"07",
		123 => x"00",
		124 => x"c1",
		125 => x"01",
		126 => x"00",
		127 => x"01",
		128 => x"81",
		129 => x"01",
		130 => x"00",
		131 => x"f4",
		132 => x"c4",
		133 => x"07",
		134 => x"c1",
		135 => x"01",
		136 => x"00",
		137 => x"01",
		138 => x"11",
		139 => x"81",
		140 => x"01",
		141 => x"00",
		142 => x"80",
		143 => x"00",
		144 => x"00",
		145 => x"00",
		146 => x"40",
		147 => x"00",
		148 => x"df",
		149 => x"01",
		150 => x"11",
		151 => x"81",
		152 => x"01",
		153 => x"05",
		154 => x"07",
		155 => x"47",
		156 => x"80",
		157 => x"c0",
		158 => x"05",
		159 => x"86",
		160 => x"a7",
		161 => x"06",
		162 => x"e8",
		163 => x"b7",
		164 => x"d8",
		165 => x"07",
		166 => x"06",
		167 => x"06",
		168 => x"e8",
		169 => x"f8",
		170 => x"00",
		171 => x"40",
		172 => x"00",
		173 => x"c1",
		174 => x"81",
		175 => x"01",
		176 => x"00",
		177 => x"01",
		178 => x"81",
		179 => x"01",
		180 => x"a4",
		181 => x"b4",
		182 => x"84",
		183 => x"c4",
		184 => x"e0",
		185 => x"f0",
		186 => x"05",
		187 => x"07",
		188 => x"47",
		189 => x"80",
		190 => x"c0",
		191 => x"05",
		192 => x"86",
		193 => x"a7",
		194 => x"06",
		195 => x"e8",
		196 => x"b7",
		197 => x"d8",
		198 => x"07",
		199 => x"06",
		200 => x"06",
		201 => x"e8",
		202 => x"f8",
		203 => x"00",
		204 => x"c1",
		205 => x"01",
		206 => x"00",
		207 => x"01",
		208 => x"11",
		209 => x"81",
		210 => x"01",
		211 => x"00",
		212 => x"df",
		213 => x"80",
		214 => x"5f",
		215 => x"00",
		216 => x"c1",
		217 => x"81",
		218 => x"01",
		219 => x"00",
		220 => x"01",
		221 => x"81",
		222 => x"01",
		223 => x"a4",
		224 => x"04",
		225 => x"80",
		226 => x"c4",
		227 => x"c4",
		228 => x"f7",
		229 => x"07",
		230 => x"09",
		231 => x"e7",
		232 => x"c4",
		233 => x"17",
		234 => x"f4",
		235 => x"c4",
		236 => x"c4",
		237 => x"f7",
		238 => x"07",
		239 => x"07",
		240 => x"00",
		241 => x"00",
		242 => x"c1",
		243 => x"01",
		244 => x"00",
		245 => x"01",
		246 => x"81",
		247 => x"01",
		248 => x"a4",
		249 => x"b4",
		250 => x"c4",
		251 => x"f4",
		252 => x"04",
		253 => x"c0",
		254 => x"c4",
		255 => x"84",
		256 => x"f7",
		257 => x"f4",
		258 => x"c4",
		259 => x"84",
		260 => x"f7",
		261 => x"f4",
		262 => x"74",
		263 => x"07",
		264 => x"f7",
		265 => x"84",
		266 => x"07",
		267 => x"87",
		268 => x"e7",
		269 => x"84",
		270 => x"17",
		271 => x"f4",
		272 => x"c4",
		273 => x"07",
		274 => x"84",
		275 => x"f7",
		276 => x"f4",
		277 => x"80",
		278 => x"84",
		279 => x"07",
		280 => x"87",
		281 => x"47",
		282 => x"09",
		283 => x"e7",
		284 => x"84",
		285 => x"f7",
		286 => x"f4",
		287 => x"84",
		288 => x"07",
		289 => x"00",
		290 => x"00",
		291 => x"c1",
		292 => x"01",
		293 => x"00",
		294 => x"01",
		295 => x"11",
		296 => x"81",
		297 => x"01",
		298 => x"df",
		299 => x"a4",
		300 => x"c4",
		301 => x"00",
		302 => x"77",
		303 => x"f7",
		304 => x"5f",
		305 => x"80",
		306 => x"80",
		307 => x"5f",
		308 => x"00",
		309 => x"c4",
		310 => x"df",
		311 => x"40",
		312 => x"1f",
		313 => x"00",
		314 => x"df",
		315 => x"00",
		316 => x"c1",
		317 => x"81",
		318 => x"01",
		319 => x"00",
		320 => x"6c",
		321 => x"77",
		322 => x"64",
		323 => x"00",
		324 => x"63",
		325 => x"00",
		326 => x"65",
		327 => x"63",
		328 => x"20",
		329 => x"75",
		330 => x"66",
		331 => x"64",
		332 => x"00",
		others => (others => '0')
	);

begin

	process(clk)
	begin
		if (rising_edge(clk)) then
			if (fetch = '1') then
				inst_out <= ram(to_integer(unsigned(addr_inst(12 downto 0))));
			end if;

			if (we = '1') then
				ram(to_integer(unsigned(addr_data(12 downto 0)))) <= data_in;
			end if;
			
			data_out <= ram(to_integer(unsigned(addr_data(12 downto 0))));
		end if;
	end process;

end behavioral ; -- arch

