library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

entity B_RAM_1 is
	port (
		clk 		: in std_logic;
		we 			: in std_logic;
		fetch		: in std_logic;
		addr_inst 	: in std_logic_vector (29 downto 0);
		addr_data	: in std_logic_vector (29 downto 0);
		data_in 	: in std_logic_vector (7 downto 0);

		inst_out 	: out std_logic_vector (7 downto 0);
		data_out 	: out std_logic_vector (7 downto 0)
	);
end B_RAM_1;

-- 8 kB BRAM
architecture behavioral of B_RAM_1 is

	type ram_type is array (0 to 8192) of std_logic_vector(7 downto 0);
	signal ram : ram_type := (
		0 => x"00",
		1 => x"80",
		2 => x"90",
		3 => x"11",
		4 => x"01",
		5 => x"00",
		6 => x"00",
		7 => x"01",
		8 => x"20",
		9 => x"00",
		10 => x"00",
		11 => x"00",
		12 => x"20",
		13 => x"01",
		14 => x"00",
		15 => x"01",
		16 => x"20",
		17 => x"22",
		18 => x"24",
		19 => x"26",
		20 => x"28",
		21 => x"2a",
		22 => x"2c",
		23 => x"2e",
		24 => x"20",
		25 => x"22",
		26 => x"24",
		27 => x"26",
		28 => x"28",
		29 => x"2a",
		30 => x"2c",
		31 => x"2e",
		32 => x"20",
		33 => x"22",
		34 => x"24",
		35 => x"26",
		36 => x"28",
		37 => x"2a",
		38 => x"2c",
		39 => x"2e",
		40 => x"20",
		41 => x"22",
		42 => x"24",
		43 => x"26",
		44 => x"28",
		45 => x"80",
		46 => x"21",
		47 => x"22",
		48 => x"22",
		49 => x"23",
		50 => x"23",
		51 => x"24",
		52 => x"24",
		53 => x"25",
		54 => x"25",
		55 => x"26",
		56 => x"26",
		57 => x"27",
		58 => x"27",
		59 => x"28",
		60 => x"28",
		61 => x"29",
		62 => x"29",
		63 => x"2a",
		64 => x"2a",
		65 => x"2b",
		66 => x"2b",
		67 => x"2c",
		68 => x"2c",
		69 => x"2d",
		70 => x"2d",
		71 => x"2e",
		72 => x"2e",
		73 => x"2f",
		74 => x"2f",
		75 => x"01",
		76 => x"80",
		77 => x"01",
		78 => x"2e",
		79 => x"04",
		80 => x"27",
		81 => x"26",
		82 => x"27",
		83 => x"85",
		84 => x"24",
		85 => x"01",
		86 => x"80",
		87 => x"01",
		88 => x"2e",
		89 => x"04",
		90 => x"26",
		91 => x"27",
		92 => x"a0",
		93 => x"00",
		94 => x"24",
		95 => x"01",
		96 => x"80",
		97 => x"01",
		98 => x"2e",
		99 => x"04",
		100 => x"26",
		101 => x"27",
		102 => x"b0",
		103 => x"00",
		104 => x"24",
		105 => x"01",
		106 => x"80",
		107 => x"01",
		108 => x"2e",
		109 => x"04",
		110 => x"26",
		111 => x"27",
		112 => x"a0",
		113 => x"00",
		114 => x"24",
		115 => x"01",
		116 => x"80",
		117 => x"01",
		118 => x"2e",
		119 => x"04",
		120 => x"26",
		121 => x"27",
		122 => x"b0",
		123 => x"00",
		124 => x"24",
		125 => x"01",
		126 => x"80",
		127 => x"01",
		128 => x"2e",
		129 => x"04",
		130 => x"27",
		131 => x"26",
		132 => x"27",
		133 => x"85",
		134 => x"24",
		135 => x"01",
		136 => x"80",
		137 => x"01",
		138 => x"26",
		139 => x"24",
		140 => x"04",
		141 => x"05",
		142 => x"00",
		143 => x"05",
		144 => x"05",
		145 => x"00",
		146 => x"00",
		147 => x"00",
		148 => x"f0",
		149 => x"01",
		150 => x"26",
		151 => x"24",
		152 => x"04",
		153 => x"07",
		154 => x"a7",
		155 => x"a7",
		156 => x"25",
		157 => x"25",
		158 => x"06",
		159 => x"88",
		160 => x"06",
		161 => x"08",
		162 => x"b8",
		163 => x"86",
		164 => x"87",
		165 => x"86",
		166 => x"07",
		167 => x"87",
		168 => x"20",
		169 => x"22",
		170 => x"05",
		171 => x"00",
		172 => x"00",
		173 => x"20",
		174 => x"24",
		175 => x"01",
		176 => x"80",
		177 => x"01",
		178 => x"2e",
		179 => x"04",
		180 => x"24",
		181 => x"26",
		182 => x"27",
		183 => x"27",
		184 => x"2c",
		185 => x"2e",
		186 => x"07",
		187 => x"a7",
		188 => x"a7",
		189 => x"25",
		190 => x"25",
		191 => x"06",
		192 => x"88",
		193 => x"06",
		194 => x"08",
		195 => x"b8",
		196 => x"86",
		197 => x"87",
		198 => x"86",
		199 => x"07",
		200 => x"87",
		201 => x"20",
		202 => x"22",
		203 => x"00",
		204 => x"24",
		205 => x"01",
		206 => x"80",
		207 => x"01",
		208 => x"26",
		209 => x"24",
		210 => x"04",
		211 => x"05",
		212 => x"f0",
		213 => x"05",
		214 => x"f0",
		215 => x"00",
		216 => x"20",
		217 => x"24",
		218 => x"01",
		219 => x"80",
		220 => x"01",
		221 => x"26",
		222 => x"04",
		223 => x"2e",
		224 => x"26",
		225 => x"00",
		226 => x"27",
		227 => x"27",
		228 => x"07",
		229 => x"c7",
		230 => x"07",
		231 => x"a0",
		232 => x"27",
		233 => x"87",
		234 => x"26",
		235 => x"27",
		236 => x"27",
		237 => x"07",
		238 => x"c7",
		239 => x"96",
		240 => x"00",
		241 => x"00",
		242 => x"24",
		243 => x"01",
		244 => x"80",
		245 => x"01",
		246 => x"26",
		247 => x"04",
		248 => x"2e",
		249 => x"2c",
		250 => x"27",
		251 => x"26",
		252 => x"24",
		253 => x"00",
		254 => x"27",
		255 => x"27",
		256 => x"77",
		257 => x"03",
		258 => x"27",
		259 => x"27",
		260 => x"57",
		261 => x"26",
		262 => x"47",
		263 => x"87",
		264 => x"f7",
		265 => x"27",
		266 => x"87",
		267 => x"87",
		268 => x"8a",
		269 => x"27",
		270 => x"87",
		271 => x"24",
		272 => x"27",
		273 => x"9a",
		274 => x"27",
		275 => x"87",
		276 => x"24",
		277 => x"00",
		278 => x"27",
		279 => x"87",
		280 => x"87",
		281 => x"c7",
		282 => x"07",
		283 => x"a0",
		284 => x"27",
		285 => x"87",
		286 => x"24",
		287 => x"27",
		288 => x"dc",
		289 => x"00",
		290 => x"00",
		291 => x"24",
		292 => x"01",
		293 => x"80",
		294 => x"01",
		295 => x"2e",
		296 => x"2c",
		297 => x"04",
		298 => x"f0",
		299 => x"26",
		300 => x"27",
		301 => x"07",
		302 => x"87",
		303 => x"16",
		304 => x"f0",
		305 => x"00",
		306 => x"05",
		307 => x"f0",
		308 => x"05",
		309 => x"25",
		310 => x"f0",
		311 => x"05",
		312 => x"f0",
		313 => x"00",
		314 => x"f0",
		315 => x"00",
		316 => x"20",
		317 => x"24",
		318 => x"01",
		319 => x"80",
		320 => x"65",
		321 => x"20",
		322 => x"6c",
		323 => x"00",
		324 => x"69",
		325 => x"0a",
		326 => x"6e",
		327 => x"65",
		328 => x"64",
		329 => x"61",
		330 => x"20",
		331 => x"6e",
		332 => x"00",
		333 => x"00",
		others => (others => '0')
	);

begin

	process(clk)
	begin
		if (rising_edge(clk)) then
			if (fetch = '1') then
				inst_out <= ram(to_integer(unsigned(addr_inst(12 downto 0))));
			end if;

			if (we = '1') then
				ram(to_integer(unsigned(addr_data(12 downto 0)))) <= data_in;
			end if;
			
			data_out <= ram(to_integer(unsigned(addr_data(12 downto 0))));
		end if;
	end process;

end behavioral ; -- arch

